module rom_meteor(
	input	[3:0]     y,
	input	[1:0]	    sprite,
	output [15:0] 	bits
);
// 16x16 Sprites (Space Meteors + Coin)
always_comb case({y, sprite})
	// 0
	6'b0000_00: bits = 16'b0000_0000_0000_0000;
	6'b0001_00: bits = 16'b0000_1111_1000_0000;
	6'b0010_00: bits = 16'b0001_1111_1110_0000;
	6'b0011_00: bits = 16'b0000_0000_1111_0000;
	6'b0100_00: bits = 16'b0010_1111_0111_1000;
	6'b0101_00: bits = 16'b0111_0111_0111_1000;
	6'b0110_00: bits = 16'b0111_1111_1001_1100;
	6'b0111_00: bits = 16'b0111_1111_1001_1100;
	6'b1000_00: bits = 16'b0111_0011_1111_1110;
	6'b1001_00: bits = 16'b0111_0111_1111_1110;
	6'b1010_00: bits = 16'b0111_1101_1111_1110;
	6'b1011_00: bits = 16'b0111_1111_1001_1100;
	6'b1100_00: bits = 16'b0011_1111_0001_1100;
	6'b1101_00: bits = 16'b0000_1111_1111_1000;
	6'b1110_00: bits = 16'b0000_0011_1111_0000;
	6'b1111_00: bits = 16'b0000_0000_0000_0000;
	//1
	6'b0000_01: bits = 16'b0000_0000_0000_0000;
	6'b0001_01: bits = 16'b0000_0111_1100_0000;
	6'b0010_01: bits = 16'b0000_1111_1110_0000;
	6'b0011_01: bits = 16'b0001_1110_1111_0000;
	6'b0100_01: bits = 16'b0011_1000_1111_1000;
	6'b0101_01: bits = 16'b0011_1001_1111_1100;
	6'b0110_01: bits = 16'b0101_1111_1110_0110;
	6'b0111_01: bits = 16'b0100_1110_1111_0110;
	6'b1000_01: bits = 16'b0111_1100_1101_1110;
	6'b1001_01: bits = 16'b0111_1111_1111_1110;
	6'b1010_01: bits = 16'b0011_1111_1111_1100;
	6'b1011_01: bits = 16'b0011_1001_1100_1000;
	6'b1100_01: bits = 16'b0000_1111_1011_0000;
	6'b1101_01: bits = 16'b0000_0111_1110_0000;
	6'b1110_01: bits = 16'b0000_0000_0000_0000;
	6'b1111_01: bits = 16'b0000_0000_0000_0000;
	//2
	6'b0000_10: bits = 16'b0000_0000_0000_0000;
	6'b0001_10: bits = 16'b0000_1111_1000_0000;
	6'b0010_10: bits = 16'b0001_1111_1110_0000;
	6'b0011_10: bits = 16'b0000_0000_1111_0000;
	6'b0100_10: bits = 16'b0010_1111_0111_1000;
	6'b0101_10: bits = 16'b0111_0111_0111_1000;
	6'b0110_10: bits = 16'b0111_1111_1001_1100;
	6'b0111_10: bits = 16'b0111_1111_1001_1100;
	6'b1000_10: bits = 16'b0011_0011_1111_1110;
	6'b1001_10: bits = 16'b0011_0111_1111_1110;
	6'b1010_10: bits = 16'b0001_1101_1111_1110;
	6'b1011_10: bits = 16'b0001_1111_1001_1100;
	6'b1100_10: bits = 16'b0000_0111_0001_1100;
	6'b1101_10: bits = 16'b0000_0011_1111_1000;
	6'b1110_10: bits = 16'b0000_0000_0111_0000;
	6'b1111_10: bits = 16'b0000_0000_0000_0000;
	//3
	6'b0000_11: bits = 16'b0000_0000_0000_0000;
	6'b0001_11: bits = 16'b0000_0000_0000_0000;
	6'b0010_11: bits = 16'b0000_0011_1000_0000;
	6'b0011_11: bits = 16'b0000_0110_1100_0000;
	6'b0100_11: bits = 16'b0000_0110_1100_0000;
	6'b0101_11: bits = 16'b0000_1100_1110_0000;
	6'b0110_11: bits = 16'b0000_1100_0110_0000;
	6'b0111_11: bits = 16'b0000_1100_0110_0000;
	6'b1000_11: bits = 16'b0000_1100_0110_0000;
	6'b1001_11: bits = 16'b0000_1100_0110_0000;
	6'b1010_11: bits = 16'b0000_1100_1110_0000;
	6'b1011_11: bits = 16'b0000_0110_1100_0000;
	6'b1100_11: bits = 16'b0000_0110_1100_0000;
	6'b1101_11: bits = 16'b0000_0011_1000_0000;
	6'b1110_11: bits = 16'b0000_0000_0000_0000;
	6'b1111_11: bits = 16'b0000_0000_0000_0000;
endcase

endmodule: rom_meteor

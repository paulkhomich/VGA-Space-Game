module rom_tail(
	input	[3:0]     y,
	input [1:0]		  frame,
	output [15:0] 	bits
);
// 16x16 Sprite (Plasma Tail from Soviet Ship)
always_comb case({frame, y})
	// frame 0
	6'b00_0000: bits = 16'b0000_0000_0000_0000;
	6'b00_0001: bits = 16'b0000_0000_0000_0000;
	6'b00_0010: bits = 16'b0000_0000_0000_0000;
	6'b00_0011: bits = 16'b0000_0000_0000_0000;
	6'b00_0100: bits = 16'b0000_0000_0000_0000;
	6'b00_0101: bits = 16'b0000_0000_0000_0111;
	6'b00_0110: bits = 16'b0000_0000_0001_1111;
	6'b00_0111: bits = 16'b0000_0000_1111_1111;
	6'b00_1000: bits = 16'b0000_0000_1111_1111;
	6'b00_1001: bits = 16'b0000_0000_0001_1111;
	6'b00_1010: bits = 16'b0000_0000_0000_0111;
	6'b00_1011: bits = 16'b0000_0000_0000_0000;
	6'b00_1100: bits = 16'b0000_0000_0000_0000;
	6'b00_1101: bits = 16'b0000_0000_0000_0000;
	6'b00_1110: bits = 16'b0000_0000_0000_0000;
	6'b00_1111: bits = 16'b0000_0000_0000_0000;
	// frame 1
	6'b01_0000: bits = 16'b0000_0000_0000_0000;
	6'b01_0001: bits = 16'b0000_0000_0000_0000;
	6'b01_0010: bits = 16'b0000_0000_0000_0000;
	6'b01_0011: bits = 16'b0000_0000_0000_0000;
	6'b01_0100: bits = 16'b0000_0000_0000_0000;
	6'b01_0101: bits = 16'b0000_0000_0000_1110;
	6'b01_0110: bits = 16'b0000_0000_0011_0000;
	6'b01_0111: bits = 16'b0000_0001_1111_1100;
	6'b01_1000: bits = 16'b0000_0001_1111_1100;
	6'b01_1001: bits = 16'b0000_0000_0011_0000;
	6'b01_1010: bits = 16'b0000_0000_0000_1110;
	6'b01_1011: bits = 16'b0000_0000_0000_0000;
	6'b01_1100: bits = 16'b0000_0000_0000_0000;
	6'b01_1101: bits = 16'b0000_0000_0000_0000;
	6'b01_1110: bits = 16'b0000_0000_0000_0000;
	6'b01_1111: bits = 16'b0000_0000_0000_0000;
	// frame 2
	6'b10_0000: bits = 16'b0000_0000_0000_0000;
	6'b10_0001: bits = 16'b0000_0000_0000_0000;
	6'b10_0010: bits = 16'b0000_0000_0000_0000;
	6'b10_0011: bits = 16'b0000_0000_0000_0000;
	6'b10_0100: bits = 16'b0000_0000_0000_0000;
	6'b10_0101: bits = 16'b0000_0000_0001_1000;
	6'b10_0110: bits = 16'b0000_0000_1111_0000;
	6'b10_0111: bits = 16'b0000_0111_1100_0001;
	6'b10_1000: bits = 16'b0000_0111_1100_0001;
	6'b10_1001: bits = 16'b0000_0000_1111_0000;
	6'b10_1010: bits = 16'b0000_0000_0001_1000;
	6'b10_1011: bits = 16'b0000_0000_0000_0000;
	6'b10_1100: bits = 16'b0000_0000_0000_0000;
	6'b10_1101: bits = 16'b0000_0000_0000_0000;
	6'b10_1110: bits = 16'b0000_0000_0000_0000;
	6'b10_1111: bits = 16'b0000_0000_0000_0000;
	// frame 3
	6'b11_0000: bits = 16'b0000_0000_0000_0000;
	6'b11_0001: bits = 16'b0000_0000_0000_0000;
	6'b11_0010: bits = 16'b0000_0000_0000_0000;
	6'b11_0011: bits = 16'b0000_0000_0000_0000;
	6'b11_0100: bits = 16'b0000_0000_0000_0000;
	6'b11_0101: bits = 16'b0000_0000_0011_0001;
	6'b11_0110: bits = 16'b0000_0001_1000_0011;
	6'b11_0111: bits = 16'b0000_0111_0001_1111;
	6'b11_1000: bits = 16'b0000_0111_0001_1111;
	6'b11_1001: bits = 16'b0000_0001_1000_0011;
	6'b11_1010: bits = 16'b0000_0000_0011_0001;
	6'b11_1011: bits = 16'b0000_0000_0000_0000;
	6'b11_1100: bits = 16'b0000_0000_0000_0000;
	6'b11_1101: bits = 16'b0000_0000_0000_0000;
	6'b11_1110: bits = 16'b0000_0000_0000_0000;
	6'b11_1111: bits = 16'b0000_0000_0000_0000;
endcase

endmodule: rom_tail

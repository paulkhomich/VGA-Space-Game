module digits(
	input [3:0]		  digit,
	input [3:0]		  line,
	output [15:0]		data_line
);	
	wire [7:0] address = {digit, line};

	always_comb 
		case (address)
			// 0
			8'b0000_0010: data_line = 16'b00111111_11111100;
			8'b0000_0011: data_line = 16'b00111111_11111100;
			8'b0000_0100: data_line = 16'b00110000_00001100;
			8'b0000_0101: data_line = 16'b00110000_00001100;
			8'b0000_0110: data_line = 16'b00110000_00001100;
			8'b0000_0111: data_line = 16'b00110000_00001100;
			8'b0000_1000: data_line = 16'b00110000_00001100;
			8'b0000_1001: data_line = 16'b00110000_00001100;
			8'b0000_1010: data_line = 16'b00110000_00001100;
			8'b0000_1011: data_line = 16'b00110000_00001100;
			8'b0000_1100: data_line = 16'b00111111_11111100;
			8'b0000_1101: data_line = 16'b00111111_11111100;
			// 1 
			8'b0001_0010: data_line = 16'b00111111_11000000;
			8'b0001_0011: data_line = 16'b00111111_11000000;
			8'b0001_0100: data_line = 16'b00000000_11000000;
			8'b0001_0101: data_line = 16'b00000000_11000000;
			8'b0001_0110: data_line = 16'b00000000_11000000;
			8'b0001_0111: data_line = 16'b00000000_11000000;
			8'b0001_1000: data_line = 16'b00000000_11000000;
			8'b0001_1001: data_line = 16'b00000000_11000000;
			8'b0001_1010: data_line = 16'b00000000_11000000;
			8'b0001_1011: data_line = 16'b00000000_11000000;
			8'b0001_1100: data_line = 16'b00111111_11111100;
			8'b0001_1101: data_line = 16'b00111111_11111100;
			// 2
			8'b0010_0010: data_line = 16'b00111111_11111100;
			8'b0010_0011: data_line = 16'b00111111_11111100;
			8'b0010_0100: data_line = 16'b00000000_00001100;
			8'b0010_0101: data_line = 16'b00000000_00001100;
			8'b0010_0110: data_line = 16'b00111111_11111100;
			8'b0010_0111: data_line = 16'b00111111_11111100;
			8'b0010_1000: data_line = 16'b00110000_00000000;
			8'b0010_1001: data_line = 16'b00110000_00000000;
			8'b0010_1010: data_line = 16'b00110000_00000000;
			8'b0010_1011: data_line = 16'b00110000_00000000;
			8'b0010_1100: data_line = 16'b00111111_11111100;
			8'b0010_1101: data_line = 16'b00111111_11111100;
			// 3
			8'b0011_0010: data_line = 16'b00111111_11111100;
			8'b0011_0011: data_line = 16'b00111111_11111100;
			8'b0011_0100: data_line = 16'b00000000_00001100;
			8'b0011_0101: data_line = 16'b00000000_00001100;
			8'b0011_0110: data_line = 16'b00111111_11111100;
			8'b0011_0111: data_line = 16'b00111111_11111100;
			8'b0011_1000: data_line = 16'b00000000_00001100;
			8'b0011_1001: data_line = 16'b00000000_00001100;
			8'b0011_1010: data_line = 16'b00000000_00001100;
			8'b0011_1011: data_line = 16'b00000000_00001100;
			8'b0011_1100: data_line = 16'b00111111_11111100;
			8'b0011_1101: data_line = 16'b00111111_11111100;
			// 4
			8'b0100_0010: data_line = 16'b00110000_00001100;
			8'b0100_0011: data_line = 16'b00110000_00001100;
			8'b0100_0100: data_line = 16'b00110000_00001100;
			8'b0100_0101: data_line = 16'b00110000_00001100;
			8'b0100_0110: data_line = 16'b00111111_11111100;
			8'b0100_0111: data_line = 16'b00111111_11111100;
			8'b0100_1000: data_line = 16'b00000000_00001100;
			8'b0100_1001: data_line = 16'b00000000_00001100;
			8'b0100_1010: data_line = 16'b00000000_00001100;
			8'b0100_1011: data_line = 16'b00000000_00001100;
			8'b0100_1100: data_line = 16'b00000000_00001100;
			8'b0100_1101: data_line = 16'b00000000_00001100;
			// 5
			8'b0101_0010: data_line = 16'b00111111_11111100;
			8'b0101_0011: data_line = 16'b00111111_11111100;
			8'b0101_0100: data_line = 16'b00110000_00000000;
			8'b0101_0101: data_line = 16'b00110000_00000000;
			8'b0101_0110: data_line = 16'b00111111_11111100;
			8'b0101_0111: data_line = 16'b00111111_11111100;
			8'b0101_1000: data_line = 16'b00000000_00001100;
			8'b0101_1001: data_line = 16'b00000000_00001100;
			8'b0101_1010: data_line = 16'b00000000_00001100;
			8'b0101_1011: data_line = 16'b00000000_00001100;
			8'b0101_1100: data_line = 16'b00111111_11111100;
			8'b0101_1101: data_line = 16'b00111111_11111100;
			// 6
			8'b0110_0010: data_line = 16'b00111111_11111100;
			8'b0110_0011: data_line = 16'b00111111_11111100;
			8'b0110_0100: data_line = 16'b00110000_00000000;
			8'b0110_0101: data_line = 16'b00110000_00000000;
			8'b0110_0110: data_line = 16'b00111111_11111100;
			8'b0110_0111: data_line = 16'b00111111_11111100;
			8'b0110_1000: data_line = 16'b00110000_00001100;
			8'b0110_1001: data_line = 16'b00110000_00001100;
			8'b0110_1010: data_line = 16'b00110000_00001100;
			8'b0110_1011: data_line = 16'b00110000_00001100;
			8'b0110_1100: data_line = 16'b00111111_11111100;
			8'b0110_1101: data_line = 16'b00111111_11111100;
			// 7
			8'b0111_0010: data_line = 16'b00111111_11111100;
			8'b0111_0011: data_line = 16'b00111111_11111100;
			8'b0111_0100: data_line = 16'b00000000_00001100;
			8'b0111_0101: data_line = 16'b00000000_00001100;
			8'b0111_0110: data_line = 16'b00000000_00001100;
			8'b0111_0111: data_line = 16'b00000000_00001100;
			8'b0111_1000: data_line = 16'b00000000_00110000;
			8'b0111_1001: data_line = 16'b00000000_00110000;
			8'b0111_1010: data_line = 16'b00000000_11000000;
			8'b0111_1011: data_line = 16'b00000000_11000000;
			8'b0111_1100: data_line = 16'b00000000_11000000;
			8'b0111_1101: data_line = 16'b00000000_11000000;
			// 8
			8'b1000_0010: data_line = 16'b00111111_11111100;
			8'b1000_0011: data_line = 16'b00111111_11111100;
			8'b1000_0100: data_line = 16'b00110000_00001100;
			8'b1000_0101: data_line = 16'b00110000_00001100;
			8'b1000_0110: data_line = 16'b00111111_11111100;
			8'b1000_0111: data_line = 16'b00111111_11111100;
			8'b1000_1000: data_line = 16'b00110000_00001100;
			8'b1000_1001: data_line = 16'b00110000_00001100;
			8'b1000_1010: data_line = 16'b00110000_00001100;
			8'b1000_1011: data_line = 16'b00110000_00001100;
			8'b1000_1100: data_line = 16'b00111111_11111100;
			8'b1000_1101: data_line = 16'b00111111_11111100;
			// 9
			8'b1001_0010: data_line = 16'b00111111_11111100;
			8'b1001_0011: data_line = 16'b00111111_11111100;
			8'b1001_0100: data_line = 16'b00110000_00001100;
			8'b1001_0101: data_line = 16'b00110000_00001100;
			8'b1001_0110: data_line = 16'b00111111_11111100;
			8'b1001_0111: data_line = 16'b00111111_11111100;
			8'b1001_1000: data_line = 16'b00000000_00001100;
			8'b1001_1001: data_line = 16'b00000000_00001100;
			8'b1001_1010: data_line = 16'b00000000_00001100;
			8'b1001_1011: data_line = 16'b00000000_00001100;
			8'b1001_1100: data_line = 16'b00111111_11111100;
			8'b1001_1101: data_line = 16'b00111111_11111100;
			// default
			default: 	 data_line = 8'b00000000_00000000;
		endcase

endmodule: digits







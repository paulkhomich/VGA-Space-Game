module rom_ship(
	input	[3:0]     y,
	output [15:0] 	bits
);
// 16x16 Sprite
// Space Ship (Soviet)
always_comb case(y)
	4'b0000: bits = 16'b0000_0000_0000_0000;
	4'b0001: bits = 16'b0000_0000_0000_0000;
	4'b0010: bits = 16'b0011_1111_1111_1100;
	4'b0011: bits = 16'b0011_1111_0000_0000;
	4'b0100: bits = 16'b0011_1000_0000_0000;
	4'b0101: bits = 16'b0111_0000_0000_0000;
	4'b0110: bits = 16'b0111_1111_0000_0000;
	4'b0111: bits = 16'b0111_1111_1111_0000;
	4'b1000: bits = 16'b0111_1111_1111_0000;
	4'b1001: bits = 16'b0111_1111_0000_0000;
	4'b1010: bits = 16'b0111_0000_0000_0000;
	4'b1011: bits = 16'b0011_1000_0000_0000;
	4'b1100: bits = 16'b0011_1111_0000_0000;
	4'b1101: bits = 16'b0011_1111_1111_1100;
	4'b1110: bits = 16'b0000_0000_0000_0000;
	4'b1111: bits = 16'b0000_0000_0000_0000;
endcase

endmodule: rom_ship
